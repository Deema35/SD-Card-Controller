module M_CRC7
(
	input wire clk,
	input wire Enable,
	input wire [47:0]  Message,
	output wire Valid,
	output reg [6:0]CRC = 'd0
);
reg [7:0] Index;
reg [7:0] Data;
reg [7:0] State = 'd0;
reg [7:0] CRC_Temp = 'd0;
reg Valid_reg = 1'b1;

assign Valid = Enable ? Valid_reg : 1'b0;


always @(posedge clk) 
begin
	if (Enable)
	begin
		if (!Valid_reg)State <= State + 1'b1;
		case(State)
			'd0: Index <= CRC_Temp ^ Message[47:40];
			'd1: CRC_Temp <= Data;
			'd2: CRC_Temp <= CRC_Temp << 1;
			'd3: Index <= CRC_Temp ^ Message[39:32];
			'd4: CRC_Temp <= Data;
			'd5: CRC_Temp <= CRC_Temp << 1;
			'd6: Index <= CRC_Temp ^ Message[31:24];
			'd7: CRC_Temp <= Data;
			'd8: CRC_Temp <= CRC_Temp << 1;
			'd9: Index <= CRC_Temp ^ Message[23:16];
			'd10: CRC_Temp <= Data;
			'd11: CRC_Temp <= CRC_Temp << 1;
			'd12: Index <= CRC_Temp ^ Message[15:8];
			'd13: 
			begin
				Valid_reg <= 1'b1;
				CRC  <= Data[6:0];
			end
		endcase
	end
	else
	begin
		State <= 1'b0;
		CRC <= 'd0;
		CRC_Temp <= 'd0;
		Valid_reg <= 1'b0;
	end
end




CRC7_ROM CRC_Table
(
	.Addr(Index),
	.data(Data)
);

endmodule

module CRC7_ROM 
#(
	parameter ADDR_WIDTH = 'd8,
	parameter DATA_WIDTH = 'd8
	
)
(   
	input wire [ADDR_WIDTH - 1:0] Addr,
	output wire [DATA_WIDTH - 1:0] data

);
 
assign data = mem[Addr];

reg [DATA_WIDTH-1:0] mem[255:0];

initial 
begin
mem[0] = 8'b00000000;
mem[1] = 8'b00001001;
mem[2] = 8'b00010010;
mem[3] = 8'b00011011;
mem[4] = 8'b00100100;
mem[5] = 8'b00101101;
mem[6] = 8'b00110110;
mem[7] = 8'b00111111;
mem[8] = 8'b01001000;
mem[9] = 8'b01000001;
mem[10] = 8'b01011010;
mem[11] = 8'b01010011;
mem[12] = 8'b01101100;
mem[13] = 8'b01100101;
mem[14] = 8'b01111110;
mem[15] = 8'b01110111;
mem[16] = 8'b00011001;
mem[17] = 8'b00010000;
mem[18] = 8'b00001011;
mem[19] = 8'b00000010;
mem[20] = 8'b00111101;
mem[21] = 8'b00110100;
mem[22] = 8'b00101111;
mem[23] = 8'b00100110;
mem[24] = 8'b01010001;
mem[25] = 8'b01011000;
mem[26] = 8'b01000011;
mem[27] = 8'b01001010;
mem[28] = 8'b01110101;
mem[29] = 8'b01111100;
mem[30] = 8'b01100111;
mem[31] = 8'b01101110;
mem[32] = 8'b00110010;
mem[33] = 8'b00111011;
mem[34] = 8'b00100000;
mem[35] = 8'b00101001;
mem[36] = 8'b00010110;
mem[37] = 8'b00011111;
mem[38] = 8'b00000100;
mem[39] = 8'b00001101;
mem[40] = 8'b01111010;
mem[41] = 8'b01110011;
mem[42] = 8'b01101000;
mem[43] = 8'b01100001;
mem[44] = 8'b01011110;
mem[45] = 8'b01010111;
mem[46] = 8'b01001100;
mem[47] = 8'b01000101;
mem[48] = 8'b00101011;
mem[49] = 8'b00100010;
mem[50] = 8'b00111001;
mem[51] = 8'b00110000;
mem[52] = 8'b00001111;
mem[53] = 8'b00000110;
mem[54] = 8'b00011101;
mem[55] = 8'b00010100;
mem[56] = 8'b01100011;
mem[57] = 8'b01101010;
mem[58] = 8'b01110001;
mem[59] = 8'b01111000;
mem[60] = 8'b01000111;
mem[61] = 8'b01001110;
mem[62] = 8'b01010101;
mem[63] = 8'b01011100;
mem[64] = 8'b01100100;
mem[65] = 8'b01101101;
mem[66] = 8'b01110110;
mem[67] = 8'b01111111;
mem[68] = 8'b01000000;
mem[69] = 8'b01001001;
mem[70] = 8'b01010010;
mem[71] = 8'b01011011;
mem[72] = 8'b00101100;
mem[73] = 8'b00100101;
mem[74] = 8'b00111110;
mem[75] = 8'b00110111;
mem[76] = 8'b00001000;
mem[77] = 8'b00000001;
mem[78] = 8'b00011010;
mem[79] = 8'b00010011;
mem[80] = 8'b01111101;
mem[81] = 8'b01110100;
mem[82] = 8'b01101111;
mem[83] = 8'b01100110;
mem[84] = 8'b01011001;
mem[85] = 8'b01010000;
mem[86] = 8'b01001011;
mem[87] = 8'b01000010;
mem[88] = 8'b00110101;
mem[89] = 8'b00111100;
mem[90] = 8'b00100111;
mem[91] = 8'b00101110;
mem[92] = 8'b00010001;
mem[93] = 8'b00011000;
mem[94] = 8'b00000011;
mem[95] = 8'b00001010;
mem[96] = 8'b01010110;
mem[97] = 8'b01011111;
mem[98] = 8'b01000100;
mem[99] = 8'b01001101;
mem[100] = 8'b01110010;
mem[101] = 8'b01111011;
mem[102] = 8'b01100000;
mem[103] = 8'b01101001;
mem[104] = 8'b00011110;
mem[105] = 8'b00010111;
mem[106] = 8'b00001100;
mem[107] = 8'b00000101;
mem[108] = 8'b00111010;
mem[109] = 8'b00110011;
mem[110] = 8'b00101000;
mem[111] = 8'b00100001;
mem[112] = 8'b01001111;
mem[113] = 8'b01000110;
mem[114] = 8'b01011101;
mem[115] = 8'b01010100;
mem[116] = 8'b01101011;
mem[117] = 8'b01100010;
mem[118] = 8'b01111001;
mem[119] = 8'b01110000;
mem[120] = 8'b00000111;
mem[121] = 8'b00001110;
mem[122] = 8'b00010101;
mem[123] = 8'b00011100;
mem[124] = 8'b00100011;
mem[125] = 8'b00101010;
mem[126] = 8'b00110001;
mem[127] = 8'b00111000;
mem[128] = 8'b01000001;
mem[129] = 8'b01001000;
mem[130] = 8'b01010011;
mem[131] = 8'b01011010;
mem[132] = 8'b01100101;
mem[133] = 8'b01101100;
mem[134] = 8'b01110111;
mem[135] = 8'b01111110;
mem[136] = 8'b00001001;
mem[137] = 8'b00000000;
mem[138] = 8'b00011011;
mem[139] = 8'b00010010;
mem[140] = 8'b00101101;
mem[141] = 8'b00100100;
mem[142] = 8'b00111111;
mem[143] = 8'b00110110;
mem[144] = 8'b01011000;
mem[145] = 8'b01010001;
mem[146] = 8'b01001010;
mem[147] = 8'b01000011;
mem[148] = 8'b01111100;
mem[149] = 8'b01110101;
mem[150] = 8'b01101110;
mem[151] = 8'b01100111;
mem[152] = 8'b00010000;
mem[153] = 8'b00011001;
mem[154] = 8'b00000010;
mem[155] = 8'b00001011;
mem[156] = 8'b00110100;
mem[157] = 8'b00111101;
mem[158] = 8'b00100110;
mem[159] = 8'b00101111;
mem[160] = 8'b01110011;
mem[161] = 8'b01111010;
mem[162] = 8'b01100001;
mem[163] = 8'b01101000;
mem[164] = 8'b01010111;
mem[165] = 8'b01011110;
mem[166] = 8'b01000101;
mem[167] = 8'b01001100;
mem[168] = 8'b00111011;
mem[169] = 8'b00110010;
mem[170] = 8'b00101001;
mem[171] = 8'b00100000;
mem[172] = 8'b00011111;
mem[173] = 8'b00010110;
mem[174] = 8'b00001101;
mem[175] = 8'b00000100;
mem[176] = 8'b01101010;
mem[177] = 8'b01100011;
mem[178] = 8'b01111000;
mem[179] = 8'b01110001;
mem[180] = 8'b01001110;
mem[181] = 8'b01000111;
mem[182] = 8'b01011100;
mem[183] = 8'b01010101;
mem[184] = 8'b00100010;
mem[185] = 8'b00101011;
mem[186] = 8'b00110000;
mem[187] = 8'b00111001;
mem[188] = 8'b00000110;
mem[189] = 8'b00001111;
mem[190] = 8'b00010100;
mem[191] = 8'b00011101;
mem[192] = 8'b00100101;
mem[193] = 8'b00101100;
mem[194] = 8'b00110111;
mem[195] = 8'b00111110;
mem[196] = 8'b00000001;
mem[197] = 8'b00001000;
mem[198] = 8'b00010011;
mem[199] = 8'b00011010;
mem[200] = 8'b01101101;
mem[201] = 8'b01100100;
mem[202] = 8'b01111111;
mem[203] = 8'b01110110;
mem[204] = 8'b01001001;
mem[205] = 8'b01000000;
mem[206] = 8'b01011011;
mem[207] = 8'b01010010;
mem[208] = 8'b00111100;
mem[209] = 8'b00110101;
mem[210] = 8'b00101110;
mem[211] = 8'b00100111;
mem[212] = 8'b00011000;
mem[213] = 8'b00010001;
mem[214] = 8'b00001010;
mem[215] = 8'b00000011;
mem[216] = 8'b01110100;
mem[217] = 8'b01111101;
mem[218] = 8'b01100110;
mem[219] = 8'b01101111;
mem[220] = 8'b01010000;
mem[221] = 8'b01011001;
mem[222] = 8'b01000010;
mem[223] = 8'b01001011;
mem[224] = 8'b00010111;
mem[225] = 8'b00011110;
mem[226] = 8'b00000101;
mem[227] = 8'b00001100;
mem[228] = 8'b00110011;
mem[229] = 8'b00111010;
mem[230] = 8'b00100001;
mem[231] = 8'b00101000;
mem[232] = 8'b01011111;
mem[233] = 8'b01010110;
mem[234] = 8'b01001101;
mem[235] = 8'b01000100;
mem[236] = 8'b01111011;
mem[237] = 8'b01110010;
mem[238] = 8'b01101001;
mem[239] = 8'b01100000;
mem[240] = 8'b00001110;
mem[241] = 8'b00000111;
mem[242] = 8'b00011100;
mem[243] = 8'b00010101;
mem[244] = 8'b00101010;
mem[245] = 8'b00100011;
mem[246] = 8'b00111000;
mem[247] = 8'b00110001;
mem[248] = 8'b01000110;
mem[249] = 8'b01001111;
mem[250] = 8'b01010100;
mem[251] = 8'b01011101;
mem[252] = 8'b01100010;
mem[253] = 8'b01101011;
mem[254] = 8'b01110000;
mem[255] = 8'b01111001;

end
endmodule