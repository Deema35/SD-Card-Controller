
module M_CRC16
#(
	DATA_STRING = 'd128
)

(
	input wire clk,
	input wire Enable,
	input wire GetData,
	input wire [7:0]  Data,
	
	output wire Valid,
	output reg [15:0]CRC = 'd0,
	
	output reg  [15:0] Index = 'd0,
	input wire [15:0] ROM_Data

);


reg [7:0] State = 'd0;
reg [15:0] CRC_Temp = 'd0;
reg Valid_reg = 1'b0;
reg [15:0]CRC_Buf = 'd0;
reg [15:0]CRC_Count = 'd0;

assign Valid = Enable ? Valid_reg : 1'b0;

localparam 	S_IDLE = 'd0,
				S_BIT_SHIFT = 'd1,
				S_INDEX_CALK = 'd2,
				S_CRC_CALK = 'd3,
				S_CRC_READY_CHECK = 'd4,
				S_COMPLITE = 'd5;
				


always @(posedge clk) 
begin
if (Enable)
	begin
		case(State)
		
		S_IDLE: if (GetData) State <= S_BIT_SHIFT;
			
			
		S_BIT_SHIFT: 
		begin
			CRC_Buf <= CRC_Temp << 8;
			CRC_Temp <= CRC_Temp >> 8;
			State <= S_INDEX_CALK;
		end
		
		S_INDEX_CALK: 
		begin
			Index <= CRC_Temp ^ Data;
			State <= S_CRC_CALK;
		end
		
		S_CRC_CALK:
		begin
			CRC_Temp <= ROM_Data ^ CRC_Buf;
			State <= S_CRC_READY_CHECK;
		end
		
		S_CRC_READY_CHECK:
		begin
			if (CRC_Count == DATA_STRING - 'd1)
			begin
				State <= S_COMPLITE;
				
				CRC  <= CRC_Temp;
			end
			else 
			begin
				State <= S_IDLE;
				CRC_Count <= CRC_Count + 1'd1;
			end
		end
		
		S_COMPLITE:
		begin
			if (Enable)
			begin
				Valid_reg <= 1'b1;
			end
			else
			begin
				Valid_reg <= 1'b0;
				State <= S_IDLE;
			end
			
		end
			
			
		endcase
	end
	else
	begin
		CRC <= 'd0;
		CRC_Temp <= 'd0;
		CRC_Buf <= 'd0;
		Valid_reg <= 1'b0;
		CRC_Count <= 1'b0;
		Index <= 'd0;
		
		State <= S_IDLE;
	end
	
end

endmodule

module M_CRC16_ROM 
#(
	parameter ADDR_WIDTH = 'd16,
	parameter DATA_WIDTH = 'd16
	
)
(   
	input wire [ADDR_WIDTH - 1:0] Index_0,
	input wire [ADDR_WIDTH - 1:0] Index_1,
	input wire [ADDR_WIDTH - 1:0] Index_2,
	input wire [ADDR_WIDTH - 1:0] Index_3,
	
	output wire [DATA_WIDTH - 1:0] ROM_Data_0,
	output wire [DATA_WIDTH - 1:0] ROM_Data_1,
	output wire [DATA_WIDTH - 1:0] ROM_Data_2,
	output wire [DATA_WIDTH - 1:0] ROM_Data_3

);
 
assign ROM_Data_0 = mem[Index_0];
assign ROM_Data_1 = mem[Index_1];
assign ROM_Data_2 = mem[Index_2];
assign ROM_Data_3 = mem[Index_3];

reg [DATA_WIDTH-1:0] mem[255:0];

initial 
begin
mem[0] = 16'b0000000000000000;
mem[1] = 16'b0001000000100001;
mem[2] = 16'b0010000001000010;
mem[3] = 16'b0011000001100011;
mem[4] = 16'b0100000010000100;
mem[5] = 16'b0101000010100101;
mem[6] = 16'b0110000011000110;
mem[7] = 16'b0111000011100111;
mem[8] = 16'b1000000100001000;
mem[9] = 16'b1001000100101001;
mem[10] = 16'b1010000101001010;
mem[11] = 16'b1011000101101011;
mem[12] = 16'b1100000110001100;
mem[13] = 16'b1101000110101101;
mem[14] = 16'b1110000111001110;
mem[15] = 16'b1111000111101111;
mem[16] = 16'b0001001000110001;
mem[17] = 16'b0000001000010000;
mem[18] = 16'b0011001001110011;
mem[19] = 16'b0010001001010010;
mem[20] = 16'b0101001010110101;
mem[21] = 16'b0100001010010100;
mem[22] = 16'b0111001011110111;
mem[23] = 16'b0110001011010110;
mem[24] = 16'b1001001100111001;
mem[25] = 16'b1000001100011000;
mem[26] = 16'b1011001101111011;
mem[27] = 16'b1010001101011010;
mem[28] = 16'b1101001110111101;
mem[29] = 16'b1100001110011100;
mem[30] = 16'b1111001111111111;
mem[31] = 16'b1110001111011110;
mem[32] = 16'b0010010001100010;
mem[33] = 16'b0011010001000011;
mem[34] = 16'b0000010000100000;
mem[35] = 16'b0001010000000001;
mem[36] = 16'b0110010011100110;
mem[37] = 16'b0111010011000111;
mem[38] = 16'b0100010010100100;
mem[39] = 16'b0101010010000101;
mem[40] = 16'b1010010101101010;
mem[41] = 16'b1011010101001011;
mem[42] = 16'b1000010100101000;
mem[43] = 16'b1001010100001001;
mem[44] = 16'b1110010111101110;
mem[45] = 16'b1111010111001111;
mem[46] = 16'b1100010110101100;
mem[47] = 16'b1101010110001101;
mem[48] = 16'b0011011001010011;
mem[49] = 16'b0010011001110010;
mem[50] = 16'b0001011000010001;
mem[51] = 16'b0000011000110000;
mem[52] = 16'b0111011011010111;
mem[53] = 16'b0110011011110110;
mem[54] = 16'b0101011010010101;
mem[55] = 16'b0100011010110100;
mem[56] = 16'b1011011101011011;
mem[57] = 16'b1010011101111010;
mem[58] = 16'b1001011100011001;
mem[59] = 16'b1000011100111000;
mem[60] = 16'b1111011111011111;
mem[61] = 16'b1110011111111110;
mem[62] = 16'b1101011110011101;
mem[63] = 16'b1100011110111100;
mem[64] = 16'b0100100011000100;
mem[65] = 16'b0101100011100101;
mem[66] = 16'b0110100010000110;
mem[67] = 16'b0111100010100111;
mem[68] = 16'b0000100001000000;
mem[69] = 16'b0001100001100001;
mem[70] = 16'b0010100000000010;
mem[71] = 16'b0011100000100011;
mem[72] = 16'b1100100111001100;
mem[73] = 16'b1101100111101101;
mem[74] = 16'b1110100110001110;
mem[75] = 16'b1111100110101111;
mem[76] = 16'b1000100101001000;
mem[77] = 16'b1001100101101001;
mem[78] = 16'b1010100100001010;
mem[79] = 16'b1011100100101011;
mem[80] = 16'b0101101011110101;
mem[81] = 16'b0100101011010100;
mem[82] = 16'b0111101010110111;
mem[83] = 16'b0110101010010110;
mem[84] = 16'b0001101001110001;
mem[85] = 16'b0000101001010000;
mem[86] = 16'b0011101000110011;
mem[87] = 16'b0010101000010010;
mem[88] = 16'b1101101111111101;
mem[89] = 16'b1100101111011100;
mem[90] = 16'b1111101110111111;
mem[91] = 16'b1110101110011110;
mem[92] = 16'b1001101101111001;
mem[93] = 16'b1000101101011000;
mem[94] = 16'b1011101100111011;
mem[95] = 16'b1010101100011010;
mem[96] = 16'b0110110010100110;
mem[97] = 16'b0111110010000111;
mem[98] = 16'b0100110011100100;
mem[99] = 16'b0101110011000101;
mem[100] = 16'b0010110000100010;
mem[101] = 16'b0011110000000011;
mem[102] = 16'b0000110001100000;
mem[103] = 16'b0001110001000001;
mem[104] = 16'b1110110110101110;
mem[105] = 16'b1111110110001111;
mem[106] = 16'b1100110111101100;
mem[107] = 16'b1101110111001101;
mem[108] = 16'b1010110100101010;
mem[109] = 16'b1011110100001011;
mem[110] = 16'b1000110101101000;
mem[111] = 16'b1001110101001001;
mem[112] = 16'b0111111010010111;
mem[113] = 16'b0110111010110110;
mem[114] = 16'b0101111011010101;
mem[115] = 16'b0100111011110100;
mem[116] = 16'b0011111000010011;
mem[117] = 16'b0010111000110010;
mem[118] = 16'b0001111001010001;
mem[119] = 16'b0000111001110000;
mem[120] = 16'b1111111110011111;
mem[121] = 16'b1110111110111110;
mem[122] = 16'b1101111111011101;
mem[123] = 16'b1100111111111100;
mem[124] = 16'b1011111100011011;
mem[125] = 16'b1010111100111010;
mem[126] = 16'b1001111101011001;
mem[127] = 16'b1000111101111000;
mem[128] = 16'b1001000110001000;
mem[129] = 16'b1000000110101001;
mem[130] = 16'b1011000111001010;
mem[131] = 16'b1010000111101011;
mem[132] = 16'b1101000100001100;
mem[133] = 16'b1100000100101101;
mem[134] = 16'b1111000101001110;
mem[135] = 16'b1110000101101111;
mem[136] = 16'b0001000010000000;
mem[137] = 16'b0000000010100001;
mem[138] = 16'b0011000011000010;
mem[139] = 16'b0010000011100011;
mem[140] = 16'b0101000000000100;
mem[141] = 16'b0100000000100101;
mem[142] = 16'b0111000001000110;
mem[143] = 16'b0110000001100111;
mem[144] = 16'b1000001110111001;
mem[145] = 16'b1001001110011000;
mem[146] = 16'b1010001111111011;
mem[147] = 16'b1011001111011010;
mem[148] = 16'b1100001100111101;
mem[149] = 16'b1101001100011100;
mem[150] = 16'b1110001101111111;
mem[151] = 16'b1111001101011110;
mem[152] = 16'b0000001010110001;
mem[153] = 16'b0001001010010000;
mem[154] = 16'b0010001011110011;
mem[155] = 16'b0011001011010010;
mem[156] = 16'b0100001000110101;
mem[157] = 16'b0101001000010100;
mem[158] = 16'b0110001001110111;
mem[159] = 16'b0111001001010110;
mem[160] = 16'b1011010111101010;
mem[161] = 16'b1010010111001011;
mem[162] = 16'b1001010110101000;
mem[163] = 16'b1000010110001001;
mem[164] = 16'b1111010101101110;
mem[165] = 16'b1110010101001111;
mem[166] = 16'b1101010100101100;
mem[167] = 16'b1100010100001101;
mem[168] = 16'b0011010011100010;
mem[169] = 16'b0010010011000011;
mem[170] = 16'b0001010010100000;
mem[171] = 16'b0000010010000001;
mem[172] = 16'b0111010001100110;
mem[173] = 16'b0110010001000111;
mem[174] = 16'b0101010000100100;
mem[175] = 16'b0100010000000101;
mem[176] = 16'b1010011111011011;
mem[177] = 16'b1011011111111010;
mem[178] = 16'b1000011110011001;
mem[179] = 16'b1001011110111000;
mem[180] = 16'b1110011101011111;
mem[181] = 16'b1111011101111110;
mem[182] = 16'b1100011100011101;
mem[183] = 16'b1101011100111100;
mem[184] = 16'b0010011011010011;
mem[185] = 16'b0011011011110010;
mem[186] = 16'b0000011010010001;
mem[187] = 16'b0001011010110000;
mem[188] = 16'b0110011001010111;
mem[189] = 16'b0111011001110110;
mem[190] = 16'b0100011000010101;
mem[191] = 16'b0101011000110100;
mem[192] = 16'b1101100101001100;
mem[193] = 16'b1100100101101101;
mem[194] = 16'b1111100100001110;
mem[195] = 16'b1110100100101111;
mem[196] = 16'b1001100111001000;
mem[197] = 16'b1000100111101001;
mem[198] = 16'b1011100110001010;
mem[199] = 16'b1010100110101011;
mem[200] = 16'b0101100001000100;
mem[201] = 16'b0100100001100101;
mem[202] = 16'b0111100000000110;
mem[203] = 16'b0110100000100111;
mem[204] = 16'b0001100011000000;
mem[205] = 16'b0000100011100001;
mem[206] = 16'b0011100010000010;
mem[207] = 16'b0010100010100011;
mem[208] = 16'b1100101101111101;
mem[209] = 16'b1101101101011100;
mem[210] = 16'b1110101100111111;
mem[211] = 16'b1111101100011110;
mem[212] = 16'b1000101111111001;
mem[213] = 16'b1001101111011000;
mem[214] = 16'b1010101110111011;
mem[215] = 16'b1011101110011010;
mem[216] = 16'b0100101001110101;
mem[217] = 16'b0101101001010100;
mem[218] = 16'b0110101000110111;
mem[219] = 16'b0111101000010110;
mem[220] = 16'b0000101011110001;
mem[221] = 16'b0001101011010000;
mem[222] = 16'b0010101010110011;
mem[223] = 16'b0011101010010010;
mem[224] = 16'b1111110100101110;
mem[225] = 16'b1110110100001111;
mem[226] = 16'b1101110101101100;
mem[227] = 16'b1100110101001101;
mem[228] = 16'b1011110110101010;
mem[229] = 16'b1010110110001011;
mem[230] = 16'b1001110111101000;
mem[231] = 16'b1000110111001001;
mem[232] = 16'b0111110000100110;
mem[233] = 16'b0110110000000111;
mem[234] = 16'b0101110001100100;
mem[235] = 16'b0100110001000101;
mem[236] = 16'b0011110010100010;
mem[237] = 16'b0010110010000011;
mem[238] = 16'b0001110011100000;
mem[239] = 16'b0000110011000001;
mem[240] = 16'b1110111100011111;
mem[241] = 16'b1111111100111110;
mem[242] = 16'b1100111101011101;
mem[243] = 16'b1101111101111100;
mem[244] = 16'b1010111110011011;
mem[245] = 16'b1011111110111010;
mem[246] = 16'b1000111111011001;
mem[247] = 16'b1001111111111000;
mem[248] = 16'b0110111000010111;
mem[249] = 16'b0111111000110110;
mem[250] = 16'b0100111001010101;
mem[251] = 16'b0101111001110100;
mem[252] = 16'b0010111010010011;
mem[253] = 16'b0011111010110010;
mem[254] = 16'b0000111011010001;
mem[255] = 16'b0001111011110000;


end

endmodule